// Copyright (c) 2022 - 2025 Advanced Micro Devices, Inc. All rights reserved.
// 
// Permission is hereby granted, free of charge, to any person obtaining a 
// copy of this software and associated documentation files (the "Software"), 
// to deal in the Software without restriction, including without limitation 
// the rights to use, copy, modify, merge, publish, distribute, sublicense, 
// and/or sell copies of the Software, and to permit persons to whom the 
// Software is furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be included in 
// all copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR 
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, 
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL 
// THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER 
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING 
// FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER 
// DEALINGS IN THE SOFTWARE.
//--------------------------------------------------------------------------

`timescale 1ps/1ps

module hw_discovery_v1_0_0_hw_discovery #(
   parameter integer C_NUM_PFS                     		     = 1,
   parameter [11:0]  C_CAP_BASE_ADDR               		     = 12'h0,
   parameter [11:0]  C_NEXT_CAP_ADDR           		         = 12'h0,
   parameter integer C_PF0_NUM_SLOTS_BAR_LAYOUT_TABLE      = 1,
   parameter integer C_PF0_BAR_INDEX               		     = 0,
   parameter [27:0]  C_PF0_LOW_OFFSET              		     = 28'h0,
   parameter [31:0]  C_PF0_HIGH_OFFSET             		     = 32'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_0                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_0                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_0                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_0           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_0           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_0            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_0                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_1                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_1                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_1                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_1           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_1           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_1            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_1                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_2                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_2                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_2                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_2           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_2           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_2            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_2                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_3                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_3                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_3                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_3           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_3           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_3            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_3                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_4                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_4                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_4                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_4           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_4           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_4            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_4                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_5                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_5                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_5                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_5           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_5           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_5            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_5                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_6                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_6                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_6                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_6           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_6           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_6            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_6                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_7                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_7                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_7                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_7           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_7           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_7            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_7                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_8                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_8                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_8                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_8           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_8           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_8            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_8                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_9                    = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_9                     = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_9                    = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_9           = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_9           = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_9            = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_9                   = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_10                   = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_10                    = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_10                   = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_10          = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_10          = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_10           = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_10                  = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_11                   = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_11                    = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_11                   = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_11          = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_11          = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_11           = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_11                  = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_12                   = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_12                    = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_12                   = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_12          = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_12          = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_12           = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_12                  = 4'h0,
   parameter [7:0]   C_PF0_ENTRY_TYPE_13                   = 8'h0,
   parameter integer C_PF0_ENTRY_BAR_13                    = 0,
   parameter [47:0]  C_PF0_ENTRY_ADDR_13                   = 48'h0,
   parameter integer C_PF0_ENTRY_MAJOR_VERSION_13          = 0,
   parameter integer C_PF0_ENTRY_MINOR_VERSION_13          = 0,
   parameter [7:0]   C_PF0_ENTRY_VERSION_TYPE_13           = 8'h0,
   parameter [3:0]   C_PF0_ENTRY_RSVD0_13                  = 4'h0,
   parameter integer C_PF0_S_AXI_ADDR_WIDTH                = 32,
   parameter integer C_PF1_NUM_SLOTS_BAR_LAYOUT_TABLE      = 1,
   parameter integer C_PF1_BAR_INDEX               		     = 0,
   parameter [27:0]  C_PF1_LOW_OFFSET              		     = 28'h0,
   parameter [31:0]  C_PF1_HIGH_OFFSET             		     = 32'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_0                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_0                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_0                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_0           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_0           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_0            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_0                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_1                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_1                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_1                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_1           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_1           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_1            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_1                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_2                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_2                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_2                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_2           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_2           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_2            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_2                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_3                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_3                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_3                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_3           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_3           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_3            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_3                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_4                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_4                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_4                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_4           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_4           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_4            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_4                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_5                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_5                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_5                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_5           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_5           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_5            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_5                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_6                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_6                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_6                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_6           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_6           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_6            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_6                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_7                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_7                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_7                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_7           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_7           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_7            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_7                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_8                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_8                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_8                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_8           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_8           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_8            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_8                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_9                    = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_9                     = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_9                    = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_9           = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_9           = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_9            = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_9                   = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_10                   = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_10                    = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_10                   = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_10          = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_10          = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_10           = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_10                  = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_11                   = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_11                    = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_11                   = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_11          = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_11          = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_11           = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_11                  = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_12                   = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_12                    = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_12                   = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_12          = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_12          = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_12           = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_12                  = 4'h0,
   parameter [7:0]   C_PF1_ENTRY_TYPE_13                   = 8'h0,
   parameter integer C_PF1_ENTRY_BAR_13                    = 0,
   parameter [47:0]  C_PF1_ENTRY_ADDR_13                   = 48'h0,
   parameter integer C_PF1_ENTRY_MAJOR_VERSION_13          = 0,
   parameter integer C_PF1_ENTRY_MINOR_VERSION_13          = 0,
   parameter [7:0]   C_PF1_ENTRY_VERSION_TYPE_13           = 8'h0,
   parameter [3:0]   C_PF1_ENTRY_RSVD0_13                  = 4'h0,
   parameter integer C_PF1_S_AXI_ADDR_WIDTH                = 32,   
   parameter integer C_PF2_NUM_SLOTS_BAR_LAYOUT_TABLE      = 1,
   parameter integer C_PF2_BAR_INDEX               		     = 0,
   parameter [27:0]  C_PF2_LOW_OFFSET              		     = 28'h0,
   parameter [31:0]  C_PF2_HIGH_OFFSET             		     = 32'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_0                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_0                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_0                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_0           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_0           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_0            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_0                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_1                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_1                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_1                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_1           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_1           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_1            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_1                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_2                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_2                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_2                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_2           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_2           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_2            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_2                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_3                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_3                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_3                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_3           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_3           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_3            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_3                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_4                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_4                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_4                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_4           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_4           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_4            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_4                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_5                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_5                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_5                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_5           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_5           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_5            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_5                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_6                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_6                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_6                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_6           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_6           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_6            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_6                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_7                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_7                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_7                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_7           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_7           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_7            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_7                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_8                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_8                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_8                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_8           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_8           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_8            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_8                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_9                    = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_9                     = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_9                    = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_9           = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_9           = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_9            = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_9                   = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_10                   = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_10                    = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_10                   = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_10          = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_10          = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_10           = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_10                  = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_11                   = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_11                    = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_11                   = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_11          = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_11          = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_11           = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_11                  = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_12                   = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_12                    = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_12                   = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_12          = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_12          = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_12           = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_12                  = 4'h0,
   parameter [7:0]   C_PF2_ENTRY_TYPE_13                   = 8'h0,
   parameter integer C_PF2_ENTRY_BAR_13                    = 0,
   parameter [47:0]  C_PF2_ENTRY_ADDR_13                   = 48'h0,
   parameter integer C_PF2_ENTRY_MAJOR_VERSION_13          = 0,
   parameter integer C_PF2_ENTRY_MINOR_VERSION_13          = 0,
   parameter [7:0]   C_PF2_ENTRY_VERSION_TYPE_13           = 8'h0,
   parameter [3:0]   C_PF2_ENTRY_RSVD0_13                  = 4'h0,
   parameter integer C_PF2_S_AXI_ADDR_WIDTH                = 32,   
   parameter integer C_PF3_NUM_SLOTS_BAR_LAYOUT_TABLE      = 1,
   parameter integer C_PF3_BAR_INDEX               		     = 0,
   parameter [27:0]  C_PF3_LOW_OFFSET              		     = 28'h0,
   parameter [31:0]  C_PF3_HIGH_OFFSET             		     = 32'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_0                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_0                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_0                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_0           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_0           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_0            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_0                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_1                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_1                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_1                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_1           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_1           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_1            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_1                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_2                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_2                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_2                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_2           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_2           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_2            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_2                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_3                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_3                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_3                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_3           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_3           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_3            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_3                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_4                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_4                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_4                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_4           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_4           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_4            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_4                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_5                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_5                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_5                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_5           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_5           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_5            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_5                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_6                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_6                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_6                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_6           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_6           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_6            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_6                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_7                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_7                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_7                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_7           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_7           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_7            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_7                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_8                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_8                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_8                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_8           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_8           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_8            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_8                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_9                    = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_9                     = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_9                    = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_9           = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_9           = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_9            = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_9                   = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_10                   = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_10                    = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_10                   = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_10          = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_10          = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_10           = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_10                  = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_11                   = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_11                    = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_11                   = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_11          = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_11          = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_11           = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_11                  = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_12                   = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_12                    = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_12                   = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_12          = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_12          = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_12           = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_12                  = 4'h0,
   parameter [7:0]   C_PF3_ENTRY_TYPE_13                   = 8'h0,
   parameter integer C_PF3_ENTRY_BAR_13                    = 0,
   parameter [47:0]  C_PF3_ENTRY_ADDR_13                   = 48'h0,
   parameter integer C_PF3_ENTRY_MAJOR_VERSION_13          = 0,
   parameter integer C_PF3_ENTRY_MINOR_VERSION_13          = 0,
   parameter [7:0]   C_PF3_ENTRY_VERSION_TYPE_13           = 8'h0,
   parameter [3:0]   C_PF3_ENTRY_RSVD0_13                  = 4'h0,
   parameter integer C_PF3_S_AXI_ADDR_WIDTH                = 32,      
   parameter         C_XDEVICEFAMILY                       = "no_family" 
   )
  (
   // Clocks & Resets
   input wire                                    aclk_pcie,
   input wire                                    aresetn_pcie,
   input wire                                    aclk_ctrl,
   input wire                                    aresetn_ctrl,
   
   // slave pcie4_cfg_ext Interface (aclk_pcie)
   input  wire [15:0]                            s_pcie4_cfg_ext_function_number,
   output wire [31:0]                            s_pcie4_cfg_ext_read_data,
   output wire                                   s_pcie4_cfg_ext_read_data_valid,
   input  wire                                   s_pcie4_cfg_ext_read_received,
   input  wire [9:0]                             s_pcie4_cfg_ext_register_number,
   input  wire [3:0]                             s_pcie4_cfg_ext_write_byte_enable,
   input  wire [31:0]                            s_pcie4_cfg_ext_write_data,
   input  wire                                   s_pcie4_cfg_ext_write_received,
   
   // slave pcie4_cfg_ext Interface (aclk_pcie)
   output wire [15:0]                            m_pcie4_cfg_ext_function_number,
   input  wire [31:0]                            m_pcie4_cfg_ext_read_data,
   input  wire                                   m_pcie4_cfg_ext_read_data_valid,
   output wire                                   m_pcie4_cfg_ext_read_received,
   output wire [9:0]                             m_pcie4_cfg_ext_register_number,
   output wire [3:0]                             m_pcie4_cfg_ext_write_byte_enable,
   output wire [31:0]                            m_pcie4_cfg_ext_write_data,
   output wire                                   m_pcie4_cfg_ext_write_received,
   
   // AXI Interface (aclk_ctrl) for PF0
   input  wire [C_PF0_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf0_awaddr,
   input  wire                                   s_axi_ctrl_pf0_awvalid,
   output wire                                   s_axi_ctrl_pf0_awready,
   input  wire [32-1:0]      s_axi_ctrl_pf0_wdata,
   input  wire [32/8-1:0]    s_axi_ctrl_pf0_wstrb,
   input  wire                                   s_axi_ctrl_pf0_wvalid,
   output wire                                   s_axi_ctrl_pf0_wready,
   output wire [1:0]                             s_axi_ctrl_pf0_bresp,
   output wire                                   s_axi_ctrl_pf0_bvalid,
   input  wire                                   s_axi_ctrl_pf0_bready,
   input  wire [C_PF0_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf0_araddr,
   input  wire                                   s_axi_ctrl_pf0_arvalid,
   output wire                                   s_axi_ctrl_pf0_arready,
   output wire [32-1:0]      s_axi_ctrl_pf0_rdata,
   output wire [1:0]                             s_axi_ctrl_pf0_rresp,
   output wire                                   s_axi_ctrl_pf0_rvalid,
   input  wire                                   s_axi_ctrl_pf0_rready,
   
   // AXI Interface (aclk_ctrl) for PF1
   input  wire [C_PF1_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf1_awaddr,
   input  wire                                   s_axi_ctrl_pf1_awvalid,
   output wire                                   s_axi_ctrl_pf1_awready,
   input  wire [32-1:0]      s_axi_ctrl_pf1_wdata,
   input  wire [32/8-1:0]    s_axi_ctrl_pf1_wstrb,
   input  wire                                   s_axi_ctrl_pf1_wvalid,
   output wire                                   s_axi_ctrl_pf1_wready,
   output wire [1:0]                             s_axi_ctrl_pf1_bresp,
   output wire                                   s_axi_ctrl_pf1_bvalid,
   input  wire                                   s_axi_ctrl_pf1_bready,
   input  wire [C_PF1_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf1_araddr,
   input  wire                                   s_axi_ctrl_pf1_arvalid,
   output wire                                   s_axi_ctrl_pf1_arready,
   output wire [32-1:0]      s_axi_ctrl_pf1_rdata,
   output wire [1:0]                             s_axi_ctrl_pf1_rresp,
   output wire                                   s_axi_ctrl_pf1_rvalid,
   input  wire                                   s_axi_ctrl_pf1_rready,
   
   // AXI Interface (aclk_ctrl) for PF2
   input  wire [C_PF2_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf2_awaddr,
   input  wire                                   s_axi_ctrl_pf2_awvalid,
   output wire                                   s_axi_ctrl_pf2_awready,
   input  wire [32-1:0]      s_axi_ctrl_pf2_wdata,
   input  wire [32/8-1:0]    s_axi_ctrl_pf2_wstrb,
   input  wire                                   s_axi_ctrl_pf2_wvalid,
   output wire                                   s_axi_ctrl_pf2_wready,
   output wire [1:0]                             s_axi_ctrl_pf2_bresp,
   output wire                                   s_axi_ctrl_pf2_bvalid,
   input  wire                                   s_axi_ctrl_pf2_bready,
   input  wire [C_PF2_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf2_araddr,
   input  wire                                   s_axi_ctrl_pf2_arvalid,
   output wire                                   s_axi_ctrl_pf2_arready,
   output wire [32-1:0]      s_axi_ctrl_pf2_rdata,
   output wire [1:0]                             s_axi_ctrl_pf2_rresp,
   output wire                                   s_axi_ctrl_pf2_rvalid,
   input  wire                                   s_axi_ctrl_pf2_rready,
   
   // AXI Interface (aclk_ctrl) for PF3
   input  wire [C_PF3_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf3_awaddr,
   input  wire                                   s_axi_ctrl_pf3_awvalid,
   output wire                                   s_axi_ctrl_pf3_awready,
   input  wire [32-1:0]      s_axi_ctrl_pf3_wdata,
   input  wire [32/8-1:0]    s_axi_ctrl_pf3_wstrb,
   input  wire                                   s_axi_ctrl_pf3_wvalid,
   output wire                                   s_axi_ctrl_pf3_wready,
   output wire [1:0]                             s_axi_ctrl_pf3_bresp,
   output wire                                   s_axi_ctrl_pf3_bvalid,
   input  wire                                   s_axi_ctrl_pf3_bready,
   input  wire [C_PF3_S_AXI_ADDR_WIDTH-1:0]      s_axi_ctrl_pf3_araddr,
   input  wire                                   s_axi_ctrl_pf3_arvalid,
   output wire                                   s_axi_ctrl_pf3_arready,
   output wire [32-1:0]      s_axi_ctrl_pf3_rdata,
   output wire [1:0]                             s_axi_ctrl_pf3_rresp,
   output wire                                   s_axi_ctrl_pf3_rvalid,
   input  wire                                   s_axi_ctrl_pf3_rready
  );
  
    hw_discovery_v1_0_0_hw_disc #(
			.C_NUM_PFS                     		    (C_NUM_PFS                     		 ),
			.C_CAP_BASE_ADDR               		    (C_CAP_BASE_ADDR               		 ),
			.C_NEXT_CAP_ADDR           		        (C_NEXT_CAP_ADDR           		     ),
			.C_PF0_NUM_SLOTS_BAR_LAYOUT_TABLE     (C_PF0_NUM_SLOTS_BAR_LAYOUT_TABLE  ),
			.C_PF0_BAR_INDEX               		    (C_PF0_BAR_INDEX               		 ),
			.C_PF0_LOW_OFFSET              		    (C_PF0_LOW_OFFSET              		 ),
			.C_PF0_HIGH_OFFSET             		    (C_PF0_HIGH_OFFSET             		 ),
			.C_PF0_ENTRY_TYPE_0                   (C_PF0_ENTRY_TYPE_0                ),
			.C_PF0_ENTRY_BAR_0                    (C_PF0_ENTRY_BAR_0                 ),
			.C_PF0_ENTRY_ADDR_0                   (C_PF0_ENTRY_ADDR_0                ),
			.C_PF0_ENTRY_MAJOR_VERSION_0          (C_PF0_ENTRY_MAJOR_VERSION_0       ),
			.C_PF0_ENTRY_MINOR_VERSION_0          (C_PF0_ENTRY_MINOR_VERSION_0       ),
			.C_PF0_ENTRY_VERSION_TYPE_0           (C_PF0_ENTRY_VERSION_TYPE_0        ),
			.C_PF0_ENTRY_RSVD0_0                  (C_PF0_ENTRY_RSVD0_0               ),
			.C_PF0_ENTRY_TYPE_1                   (C_PF0_ENTRY_TYPE_1                ),
			.C_PF0_ENTRY_BAR_1                    (C_PF0_ENTRY_BAR_1                 ),
			.C_PF0_ENTRY_ADDR_1                   (C_PF0_ENTRY_ADDR_1                ),
			.C_PF0_ENTRY_MAJOR_VERSION_1          (C_PF0_ENTRY_MAJOR_VERSION_1       ),
			.C_PF0_ENTRY_MINOR_VERSION_1          (C_PF0_ENTRY_MINOR_VERSION_1       ),
			.C_PF0_ENTRY_VERSION_TYPE_1           (C_PF0_ENTRY_VERSION_TYPE_1        ),
			.C_PF0_ENTRY_RSVD0_1                  (C_PF0_ENTRY_RSVD0_1               ),
			.C_PF0_ENTRY_TYPE_2                   (C_PF0_ENTRY_TYPE_2                ),
			.C_PF0_ENTRY_BAR_2                    (C_PF0_ENTRY_BAR_2                 ),
			.C_PF0_ENTRY_ADDR_2                   (C_PF0_ENTRY_ADDR_2                ),
			.C_PF0_ENTRY_MAJOR_VERSION_2          (C_PF0_ENTRY_MAJOR_VERSION_2       ),
			.C_PF0_ENTRY_MINOR_VERSION_2          (C_PF0_ENTRY_MINOR_VERSION_2       ),
			.C_PF0_ENTRY_VERSION_TYPE_2           (C_PF0_ENTRY_VERSION_TYPE_2        ),
			.C_PF0_ENTRY_RSVD0_2                  (C_PF0_ENTRY_RSVD0_2               ),
			.C_PF0_ENTRY_TYPE_3                   (C_PF0_ENTRY_TYPE_3                ),
			.C_PF0_ENTRY_BAR_3                    (C_PF0_ENTRY_BAR_3                 ),
			.C_PF0_ENTRY_ADDR_3                   (C_PF0_ENTRY_ADDR_3                ),
			.C_PF0_ENTRY_MAJOR_VERSION_3          (C_PF0_ENTRY_MAJOR_VERSION_3       ),
			.C_PF0_ENTRY_MINOR_VERSION_3          (C_PF0_ENTRY_MINOR_VERSION_3       ),
			.C_PF0_ENTRY_VERSION_TYPE_3           (C_PF0_ENTRY_VERSION_TYPE_3        ),
			.C_PF0_ENTRY_RSVD0_3                  (C_PF0_ENTRY_RSVD0_3               ),
			.C_PF0_ENTRY_TYPE_4                   (C_PF0_ENTRY_TYPE_4                ),
			.C_PF0_ENTRY_BAR_4                    (C_PF0_ENTRY_BAR_4                 ),
			.C_PF0_ENTRY_ADDR_4                   (C_PF0_ENTRY_ADDR_4                ),
			.C_PF0_ENTRY_MAJOR_VERSION_4          (C_PF0_ENTRY_MAJOR_VERSION_4       ),
			.C_PF0_ENTRY_MINOR_VERSION_4          (C_PF0_ENTRY_MINOR_VERSION_4       ),
			.C_PF0_ENTRY_VERSION_TYPE_4           (C_PF0_ENTRY_VERSION_TYPE_4        ),
			.C_PF0_ENTRY_RSVD0_4                  (C_PF0_ENTRY_RSVD0_4               ),
			.C_PF0_ENTRY_TYPE_5                   (C_PF0_ENTRY_TYPE_5                ),
			.C_PF0_ENTRY_BAR_5                    (C_PF0_ENTRY_BAR_5                 ),
			.C_PF0_ENTRY_ADDR_5                   (C_PF0_ENTRY_ADDR_5                ),
			.C_PF0_ENTRY_MAJOR_VERSION_5          (C_PF0_ENTRY_MAJOR_VERSION_5       ),
			.C_PF0_ENTRY_MINOR_VERSION_5          (C_PF0_ENTRY_MINOR_VERSION_5       ),
			.C_PF0_ENTRY_VERSION_TYPE_5           (C_PF0_ENTRY_VERSION_TYPE_5        ),
			.C_PF0_ENTRY_RSVD0_5                  (C_PF0_ENTRY_RSVD0_5               ),
			.C_PF0_ENTRY_TYPE_6                   (C_PF0_ENTRY_TYPE_6                ),
			.C_PF0_ENTRY_BAR_6                    (C_PF0_ENTRY_BAR_6                 ),
			.C_PF0_ENTRY_ADDR_6                   (C_PF0_ENTRY_ADDR_6                ),
			.C_PF0_ENTRY_MAJOR_VERSION_6          (C_PF0_ENTRY_MAJOR_VERSION_6       ),
			.C_PF0_ENTRY_MINOR_VERSION_6          (C_PF0_ENTRY_MINOR_VERSION_6       ),
			.C_PF0_ENTRY_VERSION_TYPE_6           (C_PF0_ENTRY_VERSION_TYPE_6        ),
			.C_PF0_ENTRY_RSVD0_6                  (C_PF0_ENTRY_RSVD0_6               ),
			.C_PF0_ENTRY_TYPE_7                   (C_PF0_ENTRY_TYPE_7                ),
			.C_PF0_ENTRY_BAR_7                    (C_PF0_ENTRY_BAR_7                 ),
			.C_PF0_ENTRY_ADDR_7                   (C_PF0_ENTRY_ADDR_7                ),
			.C_PF0_ENTRY_MAJOR_VERSION_7          (C_PF0_ENTRY_MAJOR_VERSION_7       ),
			.C_PF0_ENTRY_MINOR_VERSION_7          (C_PF0_ENTRY_MINOR_VERSION_7       ),
			.C_PF0_ENTRY_VERSION_TYPE_7           (C_PF0_ENTRY_VERSION_TYPE_7        ),
			.C_PF0_ENTRY_RSVD0_7                  (C_PF0_ENTRY_RSVD0_7               ),
			.C_PF0_ENTRY_TYPE_8                   (C_PF0_ENTRY_TYPE_8                ),
			.C_PF0_ENTRY_BAR_8                    (C_PF0_ENTRY_BAR_8                 ),
			.C_PF0_ENTRY_ADDR_8                   (C_PF0_ENTRY_ADDR_8                ),
			.C_PF0_ENTRY_MAJOR_VERSION_8          (C_PF0_ENTRY_MAJOR_VERSION_8       ),
			.C_PF0_ENTRY_MINOR_VERSION_8          (C_PF0_ENTRY_MINOR_VERSION_8       ),
			.C_PF0_ENTRY_VERSION_TYPE_8           (C_PF0_ENTRY_VERSION_TYPE_8        ),
			.C_PF0_ENTRY_RSVD0_8                  (C_PF0_ENTRY_RSVD0_8               ),
			.C_PF0_ENTRY_TYPE_9                   (C_PF0_ENTRY_TYPE_9                ),
			.C_PF0_ENTRY_BAR_9                    (C_PF0_ENTRY_BAR_9                 ),
			.C_PF0_ENTRY_ADDR_9                   (C_PF0_ENTRY_ADDR_9                ),
			.C_PF0_ENTRY_MAJOR_VERSION_9          (C_PF0_ENTRY_MAJOR_VERSION_9       ),
			.C_PF0_ENTRY_MINOR_VERSION_9          (C_PF0_ENTRY_MINOR_VERSION_9       ),
			.C_PF0_ENTRY_VERSION_TYPE_9           (C_PF0_ENTRY_VERSION_TYPE_9        ),
			.C_PF0_ENTRY_RSVD0_9                  (C_PF0_ENTRY_RSVD0_9               ),
			.C_PF0_ENTRY_TYPE_10                  (C_PF0_ENTRY_TYPE_10               ),
			.C_PF0_ENTRY_BAR_10                   (C_PF0_ENTRY_BAR_10                ),
			.C_PF0_ENTRY_ADDR_10                  (C_PF0_ENTRY_ADDR_10               ),
			.C_PF0_ENTRY_MAJOR_VERSION_10         (C_PF0_ENTRY_MAJOR_VERSION_10      ),
			.C_PF0_ENTRY_MINOR_VERSION_10         (C_PF0_ENTRY_MINOR_VERSION_10      ),
			.C_PF0_ENTRY_VERSION_TYPE_10          (C_PF0_ENTRY_VERSION_TYPE_10       ),
			.C_PF0_ENTRY_RSVD0_10                 (C_PF0_ENTRY_RSVD0_10              ),
			.C_PF0_ENTRY_TYPE_11                  (C_PF0_ENTRY_TYPE_11               ),
			.C_PF0_ENTRY_BAR_11                   (C_PF0_ENTRY_BAR_11                ),
			.C_PF0_ENTRY_ADDR_11                  (C_PF0_ENTRY_ADDR_11               ),
			.C_PF0_ENTRY_MAJOR_VERSION_11         (C_PF0_ENTRY_MAJOR_VERSION_11      ),
			.C_PF0_ENTRY_MINOR_VERSION_11         (C_PF0_ENTRY_MINOR_VERSION_11      ),
			.C_PF0_ENTRY_VERSION_TYPE_11          (C_PF0_ENTRY_VERSION_TYPE_11       ),
			.C_PF0_ENTRY_RSVD0_11                 (C_PF0_ENTRY_RSVD0_11              ),
			.C_PF0_ENTRY_TYPE_12                  (C_PF0_ENTRY_TYPE_12               ),
			.C_PF0_ENTRY_BAR_12                   (C_PF0_ENTRY_BAR_12                ),
			.C_PF0_ENTRY_ADDR_12                  (C_PF0_ENTRY_ADDR_12               ),
			.C_PF0_ENTRY_MAJOR_VERSION_12         (C_PF0_ENTRY_MAJOR_VERSION_12      ),
			.C_PF0_ENTRY_MINOR_VERSION_12         (C_PF0_ENTRY_MINOR_VERSION_12      ),
			.C_PF0_ENTRY_VERSION_TYPE_12          (C_PF0_ENTRY_VERSION_TYPE_12       ),
			.C_PF0_ENTRY_RSVD0_12                 (C_PF0_ENTRY_RSVD0_12              ),
			.C_PF0_ENTRY_TYPE_13                  (C_PF0_ENTRY_TYPE_13               ),
			.C_PF0_ENTRY_BAR_13                   (C_PF0_ENTRY_BAR_13                ),
			.C_PF0_ENTRY_ADDR_13                  (C_PF0_ENTRY_ADDR_13               ),
			.C_PF0_ENTRY_MAJOR_VERSION_13         (C_PF0_ENTRY_MAJOR_VERSION_13      ),
			.C_PF0_ENTRY_MINOR_VERSION_13         (C_PF0_ENTRY_MINOR_VERSION_13      ),
			.C_PF0_ENTRY_VERSION_TYPE_13          (C_PF0_ENTRY_VERSION_TYPE_13       ),
			.C_PF0_ENTRY_RSVD0_13                 (C_PF0_ENTRY_RSVD0_13              ),
			.C_PF0_S_AXI_ADDR_WIDTH               (C_PF0_S_AXI_ADDR_WIDTH            ),
			.C_PF1_NUM_SLOTS_BAR_LAYOUT_TABLE     (C_PF1_NUM_SLOTS_BAR_LAYOUT_TABLE  ),
			.C_PF1_BAR_INDEX               		    (C_PF1_BAR_INDEX               		 ),
			.C_PF1_LOW_OFFSET              		    (C_PF1_LOW_OFFSET              		 ),
			.C_PF1_HIGH_OFFSET             		    (C_PF1_HIGH_OFFSET             		 ),
			.C_PF1_ENTRY_TYPE_0                   (C_PF1_ENTRY_TYPE_0                ),
			.C_PF1_ENTRY_BAR_0                    (C_PF1_ENTRY_BAR_0                 ),
			.C_PF1_ENTRY_ADDR_0                   (C_PF1_ENTRY_ADDR_0                ),
			.C_PF1_ENTRY_MAJOR_VERSION_0          (C_PF1_ENTRY_MAJOR_VERSION_0       ),
			.C_PF1_ENTRY_MINOR_VERSION_0          (C_PF1_ENTRY_MINOR_VERSION_0       ),
			.C_PF1_ENTRY_VERSION_TYPE_0           (C_PF1_ENTRY_VERSION_TYPE_0        ),
			.C_PF1_ENTRY_RSVD0_0                  (C_PF1_ENTRY_RSVD0_0               ),
			.C_PF1_ENTRY_TYPE_1                   (C_PF1_ENTRY_TYPE_1                ),
			.C_PF1_ENTRY_BAR_1                    (C_PF1_ENTRY_BAR_1                 ),
			.C_PF1_ENTRY_ADDR_1                   (C_PF1_ENTRY_ADDR_1                ),
			.C_PF1_ENTRY_MAJOR_VERSION_1          (C_PF1_ENTRY_MAJOR_VERSION_1       ),
			.C_PF1_ENTRY_MINOR_VERSION_1          (C_PF1_ENTRY_MINOR_VERSION_1       ),
			.C_PF1_ENTRY_VERSION_TYPE_1           (C_PF1_ENTRY_VERSION_TYPE_1        ),
			.C_PF1_ENTRY_RSVD0_1                  (C_PF1_ENTRY_RSVD0_1               ),
			.C_PF1_ENTRY_TYPE_2                   (C_PF1_ENTRY_TYPE_2                ),
			.C_PF1_ENTRY_BAR_2                    (C_PF1_ENTRY_BAR_2                 ),
			.C_PF1_ENTRY_ADDR_2                   (C_PF1_ENTRY_ADDR_2                ),
			.C_PF1_ENTRY_MAJOR_VERSION_2          (C_PF1_ENTRY_MAJOR_VERSION_2       ),
			.C_PF1_ENTRY_MINOR_VERSION_2          (C_PF1_ENTRY_MINOR_VERSION_2       ),
			.C_PF1_ENTRY_VERSION_TYPE_2           (C_PF1_ENTRY_VERSION_TYPE_2        ),
			.C_PF1_ENTRY_RSVD0_2                  (C_PF1_ENTRY_RSVD0_2               ),
			.C_PF1_ENTRY_TYPE_3                   (C_PF1_ENTRY_TYPE_3                ),
			.C_PF1_ENTRY_BAR_3                    (C_PF1_ENTRY_BAR_3                 ),
			.C_PF1_ENTRY_ADDR_3                   (C_PF1_ENTRY_ADDR_3                ),
			.C_PF1_ENTRY_MAJOR_VERSION_3          (C_PF1_ENTRY_MAJOR_VERSION_3       ),
			.C_PF1_ENTRY_MINOR_VERSION_3          (C_PF1_ENTRY_MINOR_VERSION_3       ),
			.C_PF1_ENTRY_VERSION_TYPE_3           (C_PF1_ENTRY_VERSION_TYPE_3        ),
			.C_PF1_ENTRY_RSVD0_3                  (C_PF1_ENTRY_RSVD0_3               ),
			.C_PF1_ENTRY_TYPE_4                   (C_PF1_ENTRY_TYPE_4                ),
			.C_PF1_ENTRY_BAR_4                    (C_PF1_ENTRY_BAR_4                 ),
			.C_PF1_ENTRY_ADDR_4                   (C_PF1_ENTRY_ADDR_4                ),
			.C_PF1_ENTRY_MAJOR_VERSION_4          (C_PF1_ENTRY_MAJOR_VERSION_4       ),
			.C_PF1_ENTRY_MINOR_VERSION_4          (C_PF1_ENTRY_MINOR_VERSION_4       ),
			.C_PF1_ENTRY_VERSION_TYPE_4           (C_PF1_ENTRY_VERSION_TYPE_4        ),
			.C_PF1_ENTRY_RSVD0_4                  (C_PF1_ENTRY_RSVD0_4               ),
			.C_PF1_ENTRY_TYPE_5                   (C_PF1_ENTRY_TYPE_5                ),
			.C_PF1_ENTRY_BAR_5                    (C_PF1_ENTRY_BAR_5                 ),
			.C_PF1_ENTRY_ADDR_5                   (C_PF1_ENTRY_ADDR_5                ),
			.C_PF1_ENTRY_MAJOR_VERSION_5          (C_PF1_ENTRY_MAJOR_VERSION_5       ),
			.C_PF1_ENTRY_MINOR_VERSION_5          (C_PF1_ENTRY_MINOR_VERSION_5       ),
			.C_PF1_ENTRY_VERSION_TYPE_5           (C_PF1_ENTRY_VERSION_TYPE_5        ),
			.C_PF1_ENTRY_RSVD0_5                  (C_PF1_ENTRY_RSVD0_5               ),
			.C_PF1_ENTRY_TYPE_6                   (C_PF1_ENTRY_TYPE_6                ),
			.C_PF1_ENTRY_BAR_6                    (C_PF1_ENTRY_BAR_6                 ),
			.C_PF1_ENTRY_ADDR_6                   (C_PF1_ENTRY_ADDR_6                ),
			.C_PF1_ENTRY_MAJOR_VERSION_6          (C_PF1_ENTRY_MAJOR_VERSION_6       ),
			.C_PF1_ENTRY_MINOR_VERSION_6          (C_PF1_ENTRY_MINOR_VERSION_6       ),
			.C_PF1_ENTRY_VERSION_TYPE_6           (C_PF1_ENTRY_VERSION_TYPE_6        ),
			.C_PF1_ENTRY_RSVD0_6                  (C_PF1_ENTRY_RSVD0_6               ),
			.C_PF1_ENTRY_TYPE_7                   (C_PF1_ENTRY_TYPE_7                ),
			.C_PF1_ENTRY_BAR_7                    (C_PF1_ENTRY_BAR_7                 ),
			.C_PF1_ENTRY_ADDR_7                   (C_PF1_ENTRY_ADDR_7                ),
			.C_PF1_ENTRY_MAJOR_VERSION_7          (C_PF1_ENTRY_MAJOR_VERSION_7       ),
			.C_PF1_ENTRY_MINOR_VERSION_7          (C_PF1_ENTRY_MINOR_VERSION_7       ),
			.C_PF1_ENTRY_VERSION_TYPE_7           (C_PF1_ENTRY_VERSION_TYPE_7        ),
			.C_PF1_ENTRY_RSVD0_7                  (C_PF1_ENTRY_RSVD0_7               ),
			.C_PF1_ENTRY_TYPE_8                   (C_PF1_ENTRY_TYPE_8                ),
			.C_PF1_ENTRY_BAR_8                    (C_PF1_ENTRY_BAR_8                 ),
			.C_PF1_ENTRY_ADDR_8                   (C_PF1_ENTRY_ADDR_8                ),
			.C_PF1_ENTRY_MAJOR_VERSION_8          (C_PF1_ENTRY_MAJOR_VERSION_8       ),
			.C_PF1_ENTRY_MINOR_VERSION_8          (C_PF1_ENTRY_MINOR_VERSION_8       ),
			.C_PF1_ENTRY_VERSION_TYPE_8           (C_PF1_ENTRY_VERSION_TYPE_8        ),
			.C_PF1_ENTRY_RSVD0_8                  (C_PF1_ENTRY_RSVD0_8               ),
			.C_PF1_ENTRY_TYPE_9                   (C_PF1_ENTRY_TYPE_9                ),
			.C_PF1_ENTRY_BAR_9                    (C_PF1_ENTRY_BAR_9                 ),
			.C_PF1_ENTRY_ADDR_9                   (C_PF1_ENTRY_ADDR_9                ),
			.C_PF1_ENTRY_MAJOR_VERSION_9          (C_PF1_ENTRY_MAJOR_VERSION_9       ),
			.C_PF1_ENTRY_MINOR_VERSION_9          (C_PF1_ENTRY_MINOR_VERSION_9       ),
			.C_PF1_ENTRY_VERSION_TYPE_9           (C_PF1_ENTRY_VERSION_TYPE_9        ),
			.C_PF1_ENTRY_RSVD0_9                  (C_PF1_ENTRY_RSVD0_9               ),
			.C_PF1_ENTRY_TYPE_10                  (C_PF1_ENTRY_TYPE_10               ),
			.C_PF1_ENTRY_BAR_10                   (C_PF1_ENTRY_BAR_10                ),
			.C_PF1_ENTRY_ADDR_10                  (C_PF1_ENTRY_ADDR_10               ),
			.C_PF1_ENTRY_MAJOR_VERSION_10         (C_PF1_ENTRY_MAJOR_VERSION_10      ),
			.C_PF1_ENTRY_MINOR_VERSION_10         (C_PF1_ENTRY_MINOR_VERSION_10      ),
			.C_PF1_ENTRY_VERSION_TYPE_10          (C_PF1_ENTRY_VERSION_TYPE_10       ),
			.C_PF1_ENTRY_RSVD0_10                 (C_PF1_ENTRY_RSVD0_10              ),
			.C_PF1_ENTRY_TYPE_11                  (C_PF1_ENTRY_TYPE_11               ),
			.C_PF1_ENTRY_BAR_11                   (C_PF1_ENTRY_BAR_11                ),
			.C_PF1_ENTRY_ADDR_11                  (C_PF1_ENTRY_ADDR_11               ),
			.C_PF1_ENTRY_MAJOR_VERSION_11         (C_PF1_ENTRY_MAJOR_VERSION_11      ),
			.C_PF1_ENTRY_MINOR_VERSION_11         (C_PF1_ENTRY_MINOR_VERSION_11      ),
			.C_PF1_ENTRY_VERSION_TYPE_11          (C_PF1_ENTRY_VERSION_TYPE_11       ),
			.C_PF1_ENTRY_RSVD0_11                 (C_PF1_ENTRY_RSVD0_11              ),
			.C_PF1_ENTRY_TYPE_12                  (C_PF1_ENTRY_TYPE_12               ),
			.C_PF1_ENTRY_BAR_12                   (C_PF1_ENTRY_BAR_12                ),
			.C_PF1_ENTRY_ADDR_12                  (C_PF1_ENTRY_ADDR_12               ),
			.C_PF1_ENTRY_MAJOR_VERSION_12         (C_PF1_ENTRY_MAJOR_VERSION_12      ),
			.C_PF1_ENTRY_MINOR_VERSION_12         (C_PF1_ENTRY_MINOR_VERSION_12      ),
			.C_PF1_ENTRY_VERSION_TYPE_12          (C_PF1_ENTRY_VERSION_TYPE_12       ),
			.C_PF1_ENTRY_RSVD0_12                 (C_PF1_ENTRY_RSVD0_12              ),
			.C_PF1_ENTRY_TYPE_13                  (C_PF1_ENTRY_TYPE_13               ),
			.C_PF1_ENTRY_BAR_13                   (C_PF1_ENTRY_BAR_13                ),
			.C_PF1_ENTRY_ADDR_13                  (C_PF1_ENTRY_ADDR_13               ),
			.C_PF1_ENTRY_MAJOR_VERSION_13         (C_PF1_ENTRY_MAJOR_VERSION_13      ),
			.C_PF1_ENTRY_MINOR_VERSION_13         (C_PF1_ENTRY_MINOR_VERSION_13      ),
			.C_PF1_ENTRY_VERSION_TYPE_13          (C_PF1_ENTRY_VERSION_TYPE_13       ),
			.C_PF1_ENTRY_RSVD0_13                 (C_PF1_ENTRY_RSVD0_13              ),
			.C_PF1_S_AXI_ADDR_WIDTH               (C_PF1_S_AXI_ADDR_WIDTH            ),
			.C_PF2_NUM_SLOTS_BAR_LAYOUT_TABLE     (C_PF2_NUM_SLOTS_BAR_LAYOUT_TABLE  ),
			.C_PF2_BAR_INDEX               		    (C_PF2_BAR_INDEX               		 ),
			.C_PF2_LOW_OFFSET              		    (C_PF2_LOW_OFFSET              		 ),
			.C_PF2_HIGH_OFFSET             		    (C_PF2_HIGH_OFFSET             		 ),
			.C_PF2_ENTRY_TYPE_0                   (C_PF2_ENTRY_TYPE_0                ),
			.C_PF2_ENTRY_BAR_0                    (C_PF2_ENTRY_BAR_0                 ),
			.C_PF2_ENTRY_ADDR_0                   (C_PF2_ENTRY_ADDR_0                ),
			.C_PF2_ENTRY_MAJOR_VERSION_0          (C_PF2_ENTRY_MAJOR_VERSION_0       ),
			.C_PF2_ENTRY_MINOR_VERSION_0          (C_PF2_ENTRY_MINOR_VERSION_0       ),
			.C_PF2_ENTRY_VERSION_TYPE_0           (C_PF2_ENTRY_VERSION_TYPE_0        ),
			.C_PF2_ENTRY_RSVD0_0                  (C_PF2_ENTRY_RSVD0_0               ),
			.C_PF2_ENTRY_TYPE_1                   (C_PF2_ENTRY_TYPE_1                ),
			.C_PF2_ENTRY_BAR_1                    (C_PF2_ENTRY_BAR_1                 ),
			.C_PF2_ENTRY_ADDR_1                   (C_PF2_ENTRY_ADDR_1                ),
			.C_PF2_ENTRY_MAJOR_VERSION_1          (C_PF2_ENTRY_MAJOR_VERSION_1       ),
			.C_PF2_ENTRY_MINOR_VERSION_1          (C_PF2_ENTRY_MINOR_VERSION_1       ),
			.C_PF2_ENTRY_VERSION_TYPE_1           (C_PF2_ENTRY_VERSION_TYPE_1        ),
			.C_PF2_ENTRY_RSVD0_1                  (C_PF2_ENTRY_RSVD0_1               ),
			.C_PF2_ENTRY_TYPE_2                   (C_PF2_ENTRY_TYPE_2                ),
			.C_PF2_ENTRY_BAR_2                    (C_PF2_ENTRY_BAR_2                 ),
			.C_PF2_ENTRY_ADDR_2                   (C_PF2_ENTRY_ADDR_2                ),
			.C_PF2_ENTRY_MAJOR_VERSION_2          (C_PF2_ENTRY_MAJOR_VERSION_2       ),
			.C_PF2_ENTRY_MINOR_VERSION_2          (C_PF2_ENTRY_MINOR_VERSION_2       ),
			.C_PF2_ENTRY_VERSION_TYPE_2           (C_PF2_ENTRY_VERSION_TYPE_2        ),
			.C_PF2_ENTRY_RSVD0_2                  (C_PF2_ENTRY_RSVD0_2               ),
			.C_PF2_ENTRY_TYPE_3                   (C_PF2_ENTRY_TYPE_3                ),
			.C_PF2_ENTRY_BAR_3                    (C_PF2_ENTRY_BAR_3                 ),
			.C_PF2_ENTRY_ADDR_3                   (C_PF2_ENTRY_ADDR_3                ),
			.C_PF2_ENTRY_MAJOR_VERSION_3          (C_PF2_ENTRY_MAJOR_VERSION_3       ),
			.C_PF2_ENTRY_MINOR_VERSION_3          (C_PF2_ENTRY_MINOR_VERSION_3       ),
			.C_PF2_ENTRY_VERSION_TYPE_3           (C_PF2_ENTRY_VERSION_TYPE_3        ),
			.C_PF2_ENTRY_RSVD0_3                  (C_PF2_ENTRY_RSVD0_3               ),
			.C_PF2_ENTRY_TYPE_4                   (C_PF2_ENTRY_TYPE_4                ),
			.C_PF2_ENTRY_BAR_4                    (C_PF2_ENTRY_BAR_4                 ),
			.C_PF2_ENTRY_ADDR_4                   (C_PF2_ENTRY_ADDR_4                ),
			.C_PF2_ENTRY_MAJOR_VERSION_4          (C_PF2_ENTRY_MAJOR_VERSION_4       ),
			.C_PF2_ENTRY_MINOR_VERSION_4          (C_PF2_ENTRY_MINOR_VERSION_4       ),
			.C_PF2_ENTRY_VERSION_TYPE_4           (C_PF2_ENTRY_VERSION_TYPE_4        ),
			.C_PF2_ENTRY_RSVD0_4                  (C_PF2_ENTRY_RSVD0_4               ),
			.C_PF2_ENTRY_TYPE_5                   (C_PF2_ENTRY_TYPE_5                ),
			.C_PF2_ENTRY_BAR_5                    (C_PF2_ENTRY_BAR_5                 ),
			.C_PF2_ENTRY_ADDR_5                   (C_PF2_ENTRY_ADDR_5                ),
			.C_PF2_ENTRY_MAJOR_VERSION_5          (C_PF2_ENTRY_MAJOR_VERSION_5       ),
			.C_PF2_ENTRY_MINOR_VERSION_5          (C_PF2_ENTRY_MINOR_VERSION_5       ),
			.C_PF2_ENTRY_VERSION_TYPE_5           (C_PF2_ENTRY_VERSION_TYPE_5        ),
			.C_PF2_ENTRY_RSVD0_5                  (C_PF2_ENTRY_RSVD0_5               ),
			.C_PF2_ENTRY_TYPE_6                   (C_PF2_ENTRY_TYPE_6                ),
			.C_PF2_ENTRY_BAR_6                    (C_PF2_ENTRY_BAR_6                 ),
			.C_PF2_ENTRY_ADDR_6                   (C_PF2_ENTRY_ADDR_6                ),
			.C_PF2_ENTRY_MAJOR_VERSION_6          (C_PF2_ENTRY_MAJOR_VERSION_6       ),
			.C_PF2_ENTRY_MINOR_VERSION_6          (C_PF2_ENTRY_MINOR_VERSION_6       ),
			.C_PF2_ENTRY_VERSION_TYPE_6           (C_PF2_ENTRY_VERSION_TYPE_6        ),
			.C_PF2_ENTRY_RSVD0_6                  (C_PF2_ENTRY_RSVD0_6               ),
			.C_PF2_ENTRY_TYPE_7                   (C_PF2_ENTRY_TYPE_7                ),
			.C_PF2_ENTRY_BAR_7                    (C_PF2_ENTRY_BAR_7                 ),
			.C_PF2_ENTRY_ADDR_7                   (C_PF2_ENTRY_ADDR_7                ),
			.C_PF2_ENTRY_MAJOR_VERSION_7          (C_PF2_ENTRY_MAJOR_VERSION_7       ),
			.C_PF2_ENTRY_MINOR_VERSION_7          (C_PF2_ENTRY_MINOR_VERSION_7       ),
			.C_PF2_ENTRY_VERSION_TYPE_7           (C_PF2_ENTRY_VERSION_TYPE_7        ),
			.C_PF2_ENTRY_RSVD0_7                  (C_PF2_ENTRY_RSVD0_7               ),
			.C_PF2_ENTRY_TYPE_8                   (C_PF2_ENTRY_TYPE_8                ),
			.C_PF2_ENTRY_BAR_8                    (C_PF2_ENTRY_BAR_8                 ),
			.C_PF2_ENTRY_ADDR_8                   (C_PF2_ENTRY_ADDR_8                ),
			.C_PF2_ENTRY_MAJOR_VERSION_8          (C_PF2_ENTRY_MAJOR_VERSION_8       ),
			.C_PF2_ENTRY_MINOR_VERSION_8          (C_PF2_ENTRY_MINOR_VERSION_8       ),
			.C_PF2_ENTRY_VERSION_TYPE_8           (C_PF2_ENTRY_VERSION_TYPE_8        ),
			.C_PF2_ENTRY_RSVD0_8                  (C_PF2_ENTRY_RSVD0_8               ),
			.C_PF2_ENTRY_TYPE_9                   (C_PF2_ENTRY_TYPE_9                ),
			.C_PF2_ENTRY_BAR_9                    (C_PF2_ENTRY_BAR_9                 ),
			.C_PF2_ENTRY_ADDR_9                   (C_PF2_ENTRY_ADDR_9                ),
			.C_PF2_ENTRY_MAJOR_VERSION_9          (C_PF2_ENTRY_MAJOR_VERSION_9       ),
			.C_PF2_ENTRY_MINOR_VERSION_9          (C_PF2_ENTRY_MINOR_VERSION_9       ),
			.C_PF2_ENTRY_VERSION_TYPE_9           (C_PF2_ENTRY_VERSION_TYPE_9        ),
			.C_PF2_ENTRY_RSVD0_9                  (C_PF2_ENTRY_RSVD0_9               ),
			.C_PF2_ENTRY_TYPE_10                  (C_PF2_ENTRY_TYPE_10               ),
			.C_PF2_ENTRY_BAR_10                   (C_PF2_ENTRY_BAR_10                ),
			.C_PF2_ENTRY_ADDR_10                  (C_PF2_ENTRY_ADDR_10               ),
			.C_PF2_ENTRY_MAJOR_VERSION_10         (C_PF2_ENTRY_MAJOR_VERSION_10      ),
			.C_PF2_ENTRY_MINOR_VERSION_10         (C_PF2_ENTRY_MINOR_VERSION_10      ),
			.C_PF2_ENTRY_VERSION_TYPE_10          (C_PF2_ENTRY_VERSION_TYPE_10       ),
			.C_PF2_ENTRY_RSVD0_10                 (C_PF2_ENTRY_RSVD0_10              ),
			.C_PF2_ENTRY_TYPE_11                  (C_PF2_ENTRY_TYPE_11               ),
			.C_PF2_ENTRY_BAR_11                   (C_PF2_ENTRY_BAR_11                ),
			.C_PF2_ENTRY_ADDR_11                  (C_PF2_ENTRY_ADDR_11               ),
			.C_PF2_ENTRY_MAJOR_VERSION_11         (C_PF2_ENTRY_MAJOR_VERSION_11      ),
			.C_PF2_ENTRY_MINOR_VERSION_11         (C_PF2_ENTRY_MINOR_VERSION_11      ),
			.C_PF2_ENTRY_VERSION_TYPE_11          (C_PF2_ENTRY_VERSION_TYPE_11       ),
			.C_PF2_ENTRY_RSVD0_11                 (C_PF2_ENTRY_RSVD0_11              ),
			.C_PF2_ENTRY_TYPE_12                  (C_PF2_ENTRY_TYPE_12               ),
			.C_PF2_ENTRY_BAR_12                   (C_PF2_ENTRY_BAR_12                ),
			.C_PF2_ENTRY_ADDR_12                  (C_PF2_ENTRY_ADDR_12               ),
			.C_PF2_ENTRY_MAJOR_VERSION_12         (C_PF2_ENTRY_MAJOR_VERSION_12      ),
			.C_PF2_ENTRY_MINOR_VERSION_12         (C_PF2_ENTRY_MINOR_VERSION_12      ),
			.C_PF2_ENTRY_VERSION_TYPE_12          (C_PF2_ENTRY_VERSION_TYPE_12       ),
			.C_PF2_ENTRY_RSVD0_12                 (C_PF2_ENTRY_RSVD0_12              ),
			.C_PF2_ENTRY_TYPE_13                  (C_PF2_ENTRY_TYPE_13               ),
			.C_PF2_ENTRY_BAR_13                   (C_PF2_ENTRY_BAR_13                ),
			.C_PF2_ENTRY_ADDR_13                  (C_PF2_ENTRY_ADDR_13               ),
			.C_PF2_ENTRY_MAJOR_VERSION_13         (C_PF2_ENTRY_MAJOR_VERSION_13      ),
			.C_PF2_ENTRY_MINOR_VERSION_13         (C_PF2_ENTRY_MINOR_VERSION_13      ),
			.C_PF2_ENTRY_VERSION_TYPE_13          (C_PF2_ENTRY_VERSION_TYPE_13       ),
			.C_PF2_ENTRY_RSVD0_13                 (C_PF2_ENTRY_RSVD0_13              ),
			.C_PF2_S_AXI_ADDR_WIDTH               (C_PF2_S_AXI_ADDR_WIDTH            ),
			.C_PF3_NUM_SLOTS_BAR_LAYOUT_TABLE     (C_PF3_NUM_SLOTS_BAR_LAYOUT_TABLE  ),
			.C_PF3_BAR_INDEX               		    (C_PF3_BAR_INDEX               		 ),
			.C_PF3_LOW_OFFSET              		    (C_PF3_LOW_OFFSET              		 ),
			.C_PF3_HIGH_OFFSET             		    (C_PF3_HIGH_OFFSET             		 ),
			.C_PF3_ENTRY_TYPE_0                   (C_PF3_ENTRY_TYPE_0                ),
			.C_PF3_ENTRY_BAR_0                    (C_PF3_ENTRY_BAR_0                 ),
			.C_PF3_ENTRY_ADDR_0                   (C_PF3_ENTRY_ADDR_0                ),
			.C_PF3_ENTRY_MAJOR_VERSION_0          (C_PF3_ENTRY_MAJOR_VERSION_0       ),
			.C_PF3_ENTRY_MINOR_VERSION_0          (C_PF3_ENTRY_MINOR_VERSION_0       ),
			.C_PF3_ENTRY_VERSION_TYPE_0           (C_PF3_ENTRY_VERSION_TYPE_0        ),
			.C_PF3_ENTRY_RSVD0_0                  (C_PF3_ENTRY_RSVD0_0               ),
			.C_PF3_ENTRY_TYPE_1                   (C_PF3_ENTRY_TYPE_1                ),
			.C_PF3_ENTRY_BAR_1                    (C_PF3_ENTRY_BAR_1                 ),
			.C_PF3_ENTRY_ADDR_1                   (C_PF3_ENTRY_ADDR_1                ),
			.C_PF3_ENTRY_MAJOR_VERSION_1          (C_PF3_ENTRY_MAJOR_VERSION_1       ),
			.C_PF3_ENTRY_MINOR_VERSION_1          (C_PF3_ENTRY_MINOR_VERSION_1       ),
			.C_PF3_ENTRY_VERSION_TYPE_1           (C_PF3_ENTRY_VERSION_TYPE_1        ),
			.C_PF3_ENTRY_RSVD0_1                  (C_PF3_ENTRY_RSVD0_1               ),
			.C_PF3_ENTRY_TYPE_2                   (C_PF3_ENTRY_TYPE_2                ),
			.C_PF3_ENTRY_BAR_2                    (C_PF3_ENTRY_BAR_2                 ),
			.C_PF3_ENTRY_ADDR_2                   (C_PF3_ENTRY_ADDR_2                ),
			.C_PF3_ENTRY_MAJOR_VERSION_2          (C_PF3_ENTRY_MAJOR_VERSION_2       ),
			.C_PF3_ENTRY_MINOR_VERSION_2          (C_PF3_ENTRY_MINOR_VERSION_2       ),
			.C_PF3_ENTRY_VERSION_TYPE_2           (C_PF3_ENTRY_VERSION_TYPE_2        ),
			.C_PF3_ENTRY_RSVD0_2                  (C_PF3_ENTRY_RSVD0_2               ),
			.C_PF3_ENTRY_TYPE_3                   (C_PF3_ENTRY_TYPE_3                ),
			.C_PF3_ENTRY_BAR_3                    (C_PF3_ENTRY_BAR_3                 ),
			.C_PF3_ENTRY_ADDR_3                   (C_PF3_ENTRY_ADDR_3                ),
			.C_PF3_ENTRY_MAJOR_VERSION_3          (C_PF3_ENTRY_MAJOR_VERSION_3       ),
			.C_PF3_ENTRY_MINOR_VERSION_3          (C_PF3_ENTRY_MINOR_VERSION_3       ),
			.C_PF3_ENTRY_VERSION_TYPE_3           (C_PF3_ENTRY_VERSION_TYPE_3        ),
			.C_PF3_ENTRY_RSVD0_3                  (C_PF3_ENTRY_RSVD0_3               ),
			.C_PF3_ENTRY_TYPE_4                   (C_PF3_ENTRY_TYPE_4                ),
			.C_PF3_ENTRY_BAR_4                    (C_PF3_ENTRY_BAR_4                 ),
			.C_PF3_ENTRY_ADDR_4                   (C_PF3_ENTRY_ADDR_4                ),
			.C_PF3_ENTRY_MAJOR_VERSION_4          (C_PF3_ENTRY_MAJOR_VERSION_4       ),
			.C_PF3_ENTRY_MINOR_VERSION_4          (C_PF3_ENTRY_MINOR_VERSION_4       ),
			.C_PF3_ENTRY_VERSION_TYPE_4           (C_PF3_ENTRY_VERSION_TYPE_4        ),
			.C_PF3_ENTRY_RSVD0_4                  (C_PF3_ENTRY_RSVD0_4               ),
			.C_PF3_ENTRY_TYPE_5                   (C_PF3_ENTRY_TYPE_5                ),
			.C_PF3_ENTRY_BAR_5                    (C_PF3_ENTRY_BAR_5                 ),
			.C_PF3_ENTRY_ADDR_5                   (C_PF3_ENTRY_ADDR_5                ),
			.C_PF3_ENTRY_MAJOR_VERSION_5          (C_PF3_ENTRY_MAJOR_VERSION_5       ),
			.C_PF3_ENTRY_MINOR_VERSION_5          (C_PF3_ENTRY_MINOR_VERSION_5       ),
			.C_PF3_ENTRY_VERSION_TYPE_5           (C_PF3_ENTRY_VERSION_TYPE_5        ),
			.C_PF3_ENTRY_RSVD0_5                  (C_PF3_ENTRY_RSVD0_5               ),
			.C_PF3_ENTRY_TYPE_6                   (C_PF3_ENTRY_TYPE_6                ),
			.C_PF3_ENTRY_BAR_6                    (C_PF3_ENTRY_BAR_6                 ),
			.C_PF3_ENTRY_ADDR_6                   (C_PF3_ENTRY_ADDR_6                ),
			.C_PF3_ENTRY_MAJOR_VERSION_6          (C_PF3_ENTRY_MAJOR_VERSION_6       ),
			.C_PF3_ENTRY_MINOR_VERSION_6          (C_PF3_ENTRY_MINOR_VERSION_6       ),
			.C_PF3_ENTRY_VERSION_TYPE_6           (C_PF3_ENTRY_VERSION_TYPE_6        ),
			.C_PF3_ENTRY_RSVD0_6                  (C_PF3_ENTRY_RSVD0_6               ),
			.C_PF3_ENTRY_TYPE_7                   (C_PF3_ENTRY_TYPE_7                ),
			.C_PF3_ENTRY_BAR_7                    (C_PF3_ENTRY_BAR_7                 ),
			.C_PF3_ENTRY_ADDR_7                   (C_PF3_ENTRY_ADDR_7                ),
			.C_PF3_ENTRY_MAJOR_VERSION_7          (C_PF3_ENTRY_MAJOR_VERSION_7       ),
			.C_PF3_ENTRY_MINOR_VERSION_7          (C_PF3_ENTRY_MINOR_VERSION_7       ),
			.C_PF3_ENTRY_VERSION_TYPE_7           (C_PF3_ENTRY_VERSION_TYPE_7        ),
			.C_PF3_ENTRY_RSVD0_7                  (C_PF3_ENTRY_RSVD0_7               ),
			.C_PF3_ENTRY_TYPE_8                   (C_PF3_ENTRY_TYPE_8                ),
			.C_PF3_ENTRY_BAR_8                    (C_PF3_ENTRY_BAR_8                 ),
			.C_PF3_ENTRY_ADDR_8                   (C_PF3_ENTRY_ADDR_8                ),
			.C_PF3_ENTRY_MAJOR_VERSION_8          (C_PF3_ENTRY_MAJOR_VERSION_8       ),
			.C_PF3_ENTRY_MINOR_VERSION_8          (C_PF3_ENTRY_MINOR_VERSION_8       ),
			.C_PF3_ENTRY_VERSION_TYPE_8           (C_PF3_ENTRY_VERSION_TYPE_8        ),
			.C_PF3_ENTRY_RSVD0_8                  (C_PF3_ENTRY_RSVD0_8               ),
			.C_PF3_ENTRY_TYPE_9                   (C_PF3_ENTRY_TYPE_9                ),
			.C_PF3_ENTRY_BAR_9                    (C_PF3_ENTRY_BAR_9                 ),
			.C_PF3_ENTRY_ADDR_9                   (C_PF3_ENTRY_ADDR_9                ),
			.C_PF3_ENTRY_MAJOR_VERSION_9          (C_PF3_ENTRY_MAJOR_VERSION_9       ),
			.C_PF3_ENTRY_MINOR_VERSION_9          (C_PF3_ENTRY_MINOR_VERSION_9       ),
			.C_PF3_ENTRY_VERSION_TYPE_9           (C_PF3_ENTRY_VERSION_TYPE_9        ),
			.C_PF3_ENTRY_RSVD0_9                  (C_PF3_ENTRY_RSVD0_9               ),
			.C_PF3_ENTRY_TYPE_10                  (C_PF3_ENTRY_TYPE_10               ),
			.C_PF3_ENTRY_BAR_10                   (C_PF3_ENTRY_BAR_10                ),
			.C_PF3_ENTRY_ADDR_10                  (C_PF3_ENTRY_ADDR_10               ),
			.C_PF3_ENTRY_MAJOR_VERSION_10         (C_PF3_ENTRY_MAJOR_VERSION_10      ),
			.C_PF3_ENTRY_MINOR_VERSION_10         (C_PF3_ENTRY_MINOR_VERSION_10      ),
			.C_PF3_ENTRY_VERSION_TYPE_10          (C_PF3_ENTRY_VERSION_TYPE_10       ),
			.C_PF3_ENTRY_RSVD0_10                 (C_PF3_ENTRY_RSVD0_10              ),
			.C_PF3_ENTRY_TYPE_11                  (C_PF3_ENTRY_TYPE_11               ),
			.C_PF3_ENTRY_BAR_11                   (C_PF3_ENTRY_BAR_11                ),
			.C_PF3_ENTRY_ADDR_11                  (C_PF3_ENTRY_ADDR_11               ),
			.C_PF3_ENTRY_MAJOR_VERSION_11         (C_PF3_ENTRY_MAJOR_VERSION_11      ),
			.C_PF3_ENTRY_MINOR_VERSION_11         (C_PF3_ENTRY_MINOR_VERSION_11      ),
			.C_PF3_ENTRY_VERSION_TYPE_11          (C_PF3_ENTRY_VERSION_TYPE_11       ),
			.C_PF3_ENTRY_RSVD0_11                 (C_PF3_ENTRY_RSVD0_11              ),
			.C_PF3_ENTRY_TYPE_12                  (C_PF3_ENTRY_TYPE_12               ),
			.C_PF3_ENTRY_BAR_12                   (C_PF3_ENTRY_BAR_12                ),
			.C_PF3_ENTRY_ADDR_12                  (C_PF3_ENTRY_ADDR_12               ),
			.C_PF3_ENTRY_MAJOR_VERSION_12         (C_PF3_ENTRY_MAJOR_VERSION_12      ),
			.C_PF3_ENTRY_MINOR_VERSION_12         (C_PF3_ENTRY_MINOR_VERSION_12      ),
			.C_PF3_ENTRY_VERSION_TYPE_12          (C_PF3_ENTRY_VERSION_TYPE_12       ),
			.C_PF3_ENTRY_RSVD0_12                 (C_PF3_ENTRY_RSVD0_12              ),
			.C_PF3_ENTRY_TYPE_13                  (C_PF3_ENTRY_TYPE_13               ),
			.C_PF3_ENTRY_BAR_13                   (C_PF3_ENTRY_BAR_13                ),
			.C_PF3_ENTRY_ADDR_13                  (C_PF3_ENTRY_ADDR_13               ),
			.C_PF3_ENTRY_MAJOR_VERSION_13         (C_PF3_ENTRY_MAJOR_VERSION_13      ),
			.C_PF3_ENTRY_MINOR_VERSION_13         (C_PF3_ENTRY_MINOR_VERSION_13      ),
			.C_PF3_ENTRY_VERSION_TYPE_13          (C_PF3_ENTRY_VERSION_TYPE_13       ),
			.C_PF3_ENTRY_RSVD0_13                 (C_PF3_ENTRY_RSVD0_13              ),
			.C_PF3_S_AXI_ADDR_WIDTH               (C_PF3_S_AXI_ADDR_WIDTH            ),
			.C_XDEVICEFAMILY                      (C_XDEVICEFAMILY                   )
    ) hw_disc_inst (
      .aclk_pcie     												(aclk_pcie                         ),   
      .aresetn_pcie  												(aresetn_pcie                      ),          
      .aclk_ctrl     												(aclk_ctrl                         ),
      .aresetn_ctrl  												(aresetn_ctrl                      ),
      .s_pcie4_cfg_ext_function_number      (s_pcie4_cfg_ext_function_number   ),
      .s_pcie4_cfg_ext_read_data            (s_pcie4_cfg_ext_read_data         ),
      .s_pcie4_cfg_ext_read_data_valid      (s_pcie4_cfg_ext_read_data_valid   ),
      .s_pcie4_cfg_ext_read_received        (s_pcie4_cfg_ext_read_received     ),
      .s_pcie4_cfg_ext_register_number      (s_pcie4_cfg_ext_register_number   ),
      .s_pcie4_cfg_ext_write_byte_enable    (s_pcie4_cfg_ext_write_byte_enable ),
      .s_pcie4_cfg_ext_write_data           (s_pcie4_cfg_ext_write_data        ),
      .s_pcie4_cfg_ext_write_received       (s_pcie4_cfg_ext_write_received    ),
      .m_pcie4_cfg_ext_function_number      (m_pcie4_cfg_ext_function_number   ),
      .m_pcie4_cfg_ext_read_data            (m_pcie4_cfg_ext_read_data         ),
      .m_pcie4_cfg_ext_read_data_valid      (m_pcie4_cfg_ext_read_data_valid   ),
      .m_pcie4_cfg_ext_read_received        (m_pcie4_cfg_ext_read_received     ),
      .m_pcie4_cfg_ext_register_number      (m_pcie4_cfg_ext_register_number   ),
      .m_pcie4_cfg_ext_write_byte_enable    (m_pcie4_cfg_ext_write_byte_enable ),
      .m_pcie4_cfg_ext_write_data           (m_pcie4_cfg_ext_write_data        ),      
      .m_pcie4_cfg_ext_write_received       (m_pcie4_cfg_ext_write_received    ),
      .s_axi_ctrl_pf0_awaddr                (s_axi_ctrl_pf0_awaddr             ),
      .s_axi_ctrl_pf0_awvalid               (s_axi_ctrl_pf0_awvalid            ),
      .s_axi_ctrl_pf0_awready               (s_axi_ctrl_pf0_awready            ),
      .s_axi_ctrl_pf0_wdata                 (s_axi_ctrl_pf0_wdata              ),
      .s_axi_ctrl_pf0_wstrb                 (s_axi_ctrl_pf0_wstrb              ),
      .s_axi_ctrl_pf0_wvalid                (s_axi_ctrl_pf0_wvalid             ),
      .s_axi_ctrl_pf0_wready                (s_axi_ctrl_pf0_wready             ),
      .s_axi_ctrl_pf0_bresp                 (s_axi_ctrl_pf0_bresp              ),
      .s_axi_ctrl_pf0_bvalid                (s_axi_ctrl_pf0_bvalid             ),
      .s_axi_ctrl_pf0_bready                (s_axi_ctrl_pf0_bready             ),
      .s_axi_ctrl_pf0_araddr                (s_axi_ctrl_pf0_araddr             ),
      .s_axi_ctrl_pf0_arvalid               (s_axi_ctrl_pf0_arvalid            ),
      .s_axi_ctrl_pf0_arready               (s_axi_ctrl_pf0_arready            ),
      .s_axi_ctrl_pf0_rdata                 (s_axi_ctrl_pf0_rdata              ),
      .s_axi_ctrl_pf0_rresp                 (s_axi_ctrl_pf0_rresp              ),
      .s_axi_ctrl_pf0_rvalid                (s_axi_ctrl_pf0_rvalid             ),
      .s_axi_ctrl_pf0_rready                (s_axi_ctrl_pf0_rready             ),
      .s_axi_ctrl_pf1_awaddr                (s_axi_ctrl_pf1_awaddr             ),
      .s_axi_ctrl_pf1_awvalid               (s_axi_ctrl_pf1_awvalid            ),
      .s_axi_ctrl_pf1_awready               (s_axi_ctrl_pf1_awready            ),
      .s_axi_ctrl_pf1_wdata                 (s_axi_ctrl_pf1_wdata              ),
      .s_axi_ctrl_pf1_wstrb                 (s_axi_ctrl_pf1_wstrb              ),
      .s_axi_ctrl_pf1_wvalid                (s_axi_ctrl_pf1_wvalid             ),
      .s_axi_ctrl_pf1_wready                (s_axi_ctrl_pf1_wready             ),
      .s_axi_ctrl_pf1_bresp                 (s_axi_ctrl_pf1_bresp              ),
      .s_axi_ctrl_pf1_bvalid                (s_axi_ctrl_pf1_bvalid             ),
      .s_axi_ctrl_pf1_bready                (s_axi_ctrl_pf1_bready             ),
      .s_axi_ctrl_pf1_araddr                (s_axi_ctrl_pf1_araddr             ),
      .s_axi_ctrl_pf1_arvalid               (s_axi_ctrl_pf1_arvalid            ),
      .s_axi_ctrl_pf1_arready               (s_axi_ctrl_pf1_arready            ),
      .s_axi_ctrl_pf1_rdata                 (s_axi_ctrl_pf1_rdata              ),
      .s_axi_ctrl_pf1_rresp                 (s_axi_ctrl_pf1_rresp              ),
      .s_axi_ctrl_pf1_rvalid                (s_axi_ctrl_pf1_rvalid             ),
      .s_axi_ctrl_pf1_rready                (s_axi_ctrl_pf1_rready             ),
      .s_axi_ctrl_pf2_awaddr                (s_axi_ctrl_pf2_awaddr             ),
      .s_axi_ctrl_pf2_awvalid               (s_axi_ctrl_pf2_awvalid            ),
      .s_axi_ctrl_pf2_awready               (s_axi_ctrl_pf2_awready            ),
      .s_axi_ctrl_pf2_wdata                 (s_axi_ctrl_pf2_wdata              ),
      .s_axi_ctrl_pf2_wstrb                 (s_axi_ctrl_pf2_wstrb              ),
      .s_axi_ctrl_pf2_wvalid                (s_axi_ctrl_pf2_wvalid             ),
      .s_axi_ctrl_pf2_wready                (s_axi_ctrl_pf2_wready             ),
      .s_axi_ctrl_pf2_bresp                 (s_axi_ctrl_pf2_bresp              ),
      .s_axi_ctrl_pf2_bvalid                (s_axi_ctrl_pf2_bvalid             ),
      .s_axi_ctrl_pf2_bready                (s_axi_ctrl_pf2_bready             ),
      .s_axi_ctrl_pf2_araddr                (s_axi_ctrl_pf2_araddr             ),
      .s_axi_ctrl_pf2_arvalid               (s_axi_ctrl_pf2_arvalid            ),
      .s_axi_ctrl_pf2_arready               (s_axi_ctrl_pf2_arready            ),
      .s_axi_ctrl_pf2_rdata                 (s_axi_ctrl_pf2_rdata              ),
      .s_axi_ctrl_pf2_rresp                 (s_axi_ctrl_pf2_rresp              ),
      .s_axi_ctrl_pf2_rvalid                (s_axi_ctrl_pf2_rvalid             ),
      .s_axi_ctrl_pf2_rready                (s_axi_ctrl_pf2_rready             ),
      .s_axi_ctrl_pf3_awaddr                (s_axi_ctrl_pf3_awaddr             ),
      .s_axi_ctrl_pf3_awvalid               (s_axi_ctrl_pf3_awvalid            ),
      .s_axi_ctrl_pf3_awready               (s_axi_ctrl_pf3_awready            ),
      .s_axi_ctrl_pf3_wdata                 (s_axi_ctrl_pf3_wdata              ),
      .s_axi_ctrl_pf3_wstrb                 (s_axi_ctrl_pf3_wstrb              ),
      .s_axi_ctrl_pf3_wvalid                (s_axi_ctrl_pf3_wvalid             ),
      .s_axi_ctrl_pf3_wready                (s_axi_ctrl_pf3_wready             ),
      .s_axi_ctrl_pf3_bresp                 (s_axi_ctrl_pf3_bresp              ),
      .s_axi_ctrl_pf3_bvalid                (s_axi_ctrl_pf3_bvalid             ),
      .s_axi_ctrl_pf3_bready                (s_axi_ctrl_pf3_bready             ),
      .s_axi_ctrl_pf3_araddr                (s_axi_ctrl_pf3_araddr             ),
      .s_axi_ctrl_pf3_arvalid               (s_axi_ctrl_pf3_arvalid            ),
      .s_axi_ctrl_pf3_arready               (s_axi_ctrl_pf3_arready            ),
      .s_axi_ctrl_pf3_rdata                 (s_axi_ctrl_pf3_rdata              ),
      .s_axi_ctrl_pf3_rresp                 (s_axi_ctrl_pf3_rresp              ),
      .s_axi_ctrl_pf3_rvalid                (s_axi_ctrl_pf3_rvalid             ),
      .s_axi_ctrl_pf3_rready                (s_axi_ctrl_pf3_rready             )
    );
    
endmodule
